module Instruction_Memory (A , 
            RD );

/********************** parameters **********************/

/********************** input declaration **********************/
input wire [31 : 0] A;

/********************** output declaration **********************/
output wire [31 : 0] RD;

/********************** Memory Declaration **********************/
reg [31:0] DATA [255:0]; 

/**********************   descriptin   **********************/
assign RD = DATA[A[9:2]];

initial 
begin
    DATA[0]  = 32'b00000000101000000000000010010011;  // addi x1, x0, 10
    DATA[1]  = 32'b00000001010000000000000100010011;  // addi x2, x0, 20
    DATA[2]  = 32'b00000010100000000000000110010011;  // addi x3, x0, 40
    DATA[3]  = 32'b00000101000000000000001000010011;  // addi x4, x0, 80
    DATA[4]  = 32'b00001010000000000000001010010011;  // addi x5, x0, 160
    DATA[5]  = 32'b00000000000100000010000000100011;  // sw x1, 0(x0)
    DATA[6]  = 32'b00000000001000000010001000100011;  // sw x2, 4(x0)
    DATA[7]  = 32'b00000000001100000010010000100011;  // sw x3, 8(x0)
    DATA[8]  = 32'b00000000010000000010011000100011;  // sw x4, 12(x0)
    DATA[9]  = 32'b00000000010100000010011000100011;  // sw x5, 12(x0)
    DATA[10] = 32'b00000000000000000010010100000011;  // lw x10, 0(x0)
    DATA[11] = 32'b00000000010000000010010110000011;  // lw x11, 4(x0)
    DATA[12] = 32'b00000000100000000010011000000011;  // lw x12, 8(x0)
    DATA[13] = 32'b00000000110000000010011010000011;  // lw x13, 12(x0)
    DATA[14] = 32'b00000000010000000010011000100011;  // sw x4, 12(x0)
    /*
    DATA[0]  = 32'h0050_0113;
    DATA[1]  = 32'h00C0_0193;
    DATA[2]  = 32'hFF71_8393;
    DATA[3]  = 32'h0023_E233;
    DATA[4]  = 32'h0041_F2B3;
    DATA[5]  = 32'h0042_82B3;
    DATA[6]  = 32'h0272_8863;
    DATA[7]  = 32'h0041_A233;
    DATA[8]  = 32'h0002_0463;
    DATA[9]  = 32'h0000_0293;
    DATA[10] = 32'h0023_A233;
    DATA[11] = 32'h0052_03B3;
    DATA[12] = 32'h4023_83B3;
    DATA[13] = 32'h0471_AA23;
    DATA[14] = 32'h0600_2103;
    DATA[15] = 32'h0051_04B3;
    DATA[16] = 32'h0080_01EF;
    DATA[17] = 32'h0010_0113;
    DATA[18] = 32'h0091_0133;
    DATA[19] = 32'h0221_A023;
    DATA[20] = 32'h0021_0063;*/

    /*
    main: addi x2, x0, 5 # x2 = 5 0 00500113
        addi x3, x0, 12 # x3 = 12 4 00C00193
        addi x7, x3, -9 # x7 = (12 - 9) = 3 8 FF718393
        or x4, x7, x2 # x4 = (3 OR 5) = 7 C 0023E233
        and x5, x3, x4 # x5 = (12 AND 7) = 4 10 0041F2B3
        add x5, x5, x4 # x5 = 4 + 7 = 11 14 004282B3
        beq x5, x7, end # shouldn't be taken 18 02728863
        slt x4, x3, x4 # x4 = (12 < 7) = 0 1C 0041A233
        beq x4, x0, around # should be taken 20 00020463
        addi x5, x0, 0 # shouldn't execute 24 00000293
    around: slt x4, x7, x2 # x4 = (3 < 5) = 1 28 0023A233
        add x7, x4, x5 # x7 = (1 + 11) = 12 2C 005203B3
        sub x7, x7, x2 # x7 = (12 - 5) = 7 30 402383B3
        sw x7, 84(x3) # [96] = 7 34 0471AA23
        lw x2, 96(x0) # x2 = [96] = 7 38 06002103
        add x9, x2, x5 # x9 = (7 + 11) = 18 3C 005104B3
        jal x3, end # jump to end, x3 = 0x44 40 008001EF
        addi x2, x0, 1 # shouldn't execute 44 00100113
    end: add x2, x2, x9 # x2 = (7 + 18) = 25 48 4C    00910133
         sw x2, 0x20(x3) # [100] = 25 0221A023
    done: beq x2, x2, done # infinite loop 50 00210063
    */
end

endmodule
